*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_OTA_lpe.spi
#else
.include ../../../work/xsch/CNR_OTA.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  0  dc {AVDD}


vlp1 lpci lpco dc 0

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

.include ../load.spi


.include ../../../../cpdk/ngspice/balun.spi
xb1 LPO VCM VOP VON balun
xb2 LPI VCM LOP LON balun


.include ../../../../cpdk/ngspice/tian_subckt.lib
X999 LPI LPO loopgainprobe

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

.save v(xdut.vbn1) v(xdut.vbn2) v(xdut.vbn) v(xdut.vcn)
.save v(xdut.vbp1) v(xdut.vbp2) v(xdut.vbp) v(xdut.vcp)
.save v(xdut.vconp) v(xdut.vconn) v(xdut.vcopn) v(xdut.vcopp)
.save v(xdut.vs)
.save v(xdut.vcbp)
.save v(xdut.vco) v(xdut.vcref)
.save v(xdut.vcs)
.save v(von) v(vop) v(vin) v(vip) v(ibpsr_5u) v(vdd_1v8) v(vss) v(vsin) v(vsip)

.save V(X999.x) I(v.X999.Vi)
.save v(LPO) v(LPI) v(LOP) V(LON)
.save v(AVDD)
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100n 4u 0
op
write {cicname}_op.raw

*----------------------------------------------------------------
* LSTB analysis
*----------------------------------------------------------------
* Set voltage AC to 1
ac dec 50 1 0.1G

* Set Current to 1
alter i.X999.Ii acmag=1
alter v.X999.Vi acmag=0
ac dec 50 1 0.1G

let lg_mag = db(tian_loop())
let lg_phase = 180*cph(tian_loop())/pi


write

quit

.endc

.end
